module geofence ( clk,reset,X,Y,valid,is_inside);
input clk;
input reset;
input [9:0] X;
input [9:0] Y;
output valid;
output is_inside;
//reg valid;
//reg is_inside;

always @(posedge clk or posedge reset) begin

end

always @(posedge clk or posedge reset) begin
%{}
end

always @(posedge clk or posedge reset) begin
${}
end

always @(posedge clk or posedge reset) begin

end

always @(posedge clk or posedge reset) begin
    
end

if()begin

end
else begin
end

if()begin

end
else begin

end
endmodule

