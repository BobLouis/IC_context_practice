`timescale 1ns/10ps
module CS(Y, X, reset, clk);

    input clk, reset; 
    input 	[7:0] X;
    output reg	[9:0] Y;
    reg 

endmodule