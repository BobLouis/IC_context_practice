module triangle (clk, reset, nt, xi, yi, busy, po, xo, yo);
   input clk, reset, nt;
   input [2:0] xi, yi;
   output busy, po;
   output [2:0] xo, yo;
  

   
endmodule